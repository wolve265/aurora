`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 08.02.2023 20:15:32
// Design Name:
// Module Name: pseudo_random_integer_generator
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module pseudo_random_integer_generator(
    input logic clk,
    output logic pseudo_random_bit,
    output logic [7:0] pseudo_random_integer
    );

    // TODO: implement pseudo_random

endmodule
